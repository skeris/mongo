module bson

