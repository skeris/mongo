module description

struct SelectedServer {
	
}